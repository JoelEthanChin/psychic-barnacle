module fsm(x, y, z);

  
